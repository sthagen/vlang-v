module fasthttp

import net

#include <sys/epoll.h>
#include <sys/sendfile.h>
#include <sys/stat.h>
#include <netinet/tcp.h>

fn C.accept4(sockfd i32, addr &net.Addr, addrlen &u32, flags i32) i32

fn C.epoll_create1(__flags i32) i32

fn C.epoll_ctl(__epfd i32, __op i32, __fd i32, __event &C.epoll_event) i32

fn C.epoll_wait(__epfd i32, __events &C.epoll_event, __maxevents i32, __timeout i32) i32

fn C.sendfile(out_fd i32, in_fd i32, offset &i64, count usize) i32

fn C.fstat(fd i32, buf &C.stat) i32

@[typedef]
union C.epoll_data_t {
	ptr voidptr
	fd  int
	u32 u32
	u64 u64
}

struct C.epoll_event {
	events u32
	data   C.epoll_data_t
}

struct Server {
pub:
	family                  net.AddrFamily = .ip6
	port                    int            = 3000
	max_request_buffer_size int            = 8192
	user_data               voidptr
mut:
	listen_fds      []int    = []int{len: max_thread_pool_size, cap: max_thread_pool_size}
	epoll_fds       []int    = []int{len: max_thread_pool_size, cap: max_thread_pool_size}
	threads         []thread = []thread{len: max_thread_pool_size, cap: max_thread_pool_size}
	request_handler fn (HttpRequest) !HttpResponse @[required]
}

// new_server creates and initializes a new Server instance.
pub fn new_server(config ServerConfig) !&Server {
	if config.max_request_buffer_size <= 0 {
		return error('max_request_buffer_size must be greater than 0')
	}
	mut server := &Server{
		family:                  config.family
		port:                    config.port
		max_request_buffer_size: config.max_request_buffer_size
		user_data:               config.user_data
		request_handler:         config.handler
	}
	unsafe {
		server.listen_fds.flags.set(.noslices | .noshrink | .nogrow)
		server.epoll_fds.flags.set(.noslices | .noshrink | .nogrow)
		server.threads.flags.set(.noslices | .noshrink | .nogrow)
	}
	return server
}

fn set_blocking(fd int, blocking bool) {
	flags := C.fcntl(fd, C.F_GETFL, 0)
	if flags == -1 {
		// TODO: better error handling
		eprintln(@LOCATION)
		return
	}
	if blocking {
		// This removes the O_NONBLOCK flag from flags and set it.
		C.fcntl(fd, C.F_SETFL, flags & ~C.O_NONBLOCK)
	} else {
		// This adds the O_NONBLOCK flag from flags and set it.
		C.fcntl(fd, C.F_SETFL, flags | C.O_NONBLOCK)
	}
}

fn close_socket(fd int) bool {
	ret := C.close(fd)
	if ret == -1 {
		if C.errno == C.EINTR {
			// Interrupted by signal, retry is safe
			return close_socket(fd)
		}
		eprintln('ERROR: close(fd=${fd}) failed with errno=${C.errno}')
		return false
	}
	return true
}

fn create_server_socket(server Server) int {
	// Create a socket with non-blocking mode
	server_fd := C.socket(server.family, net.SocketType.tcp, 0)
	if server_fd < 0 {
		eprintln(@LOCATION)
		C.perror(c'Socket creation failed')
		return -1
	}

	set_blocking(server_fd, false)

	// Enable SO_REUSEADDR and SO_REUSEPORT
	opt := 1
	if C.setsockopt(server_fd, C.SOL_SOCKET, C.SO_REUSEADDR, &opt, sizeof(opt)) < 0 {
		eprintln(@LOCATION)
		C.perror(c'setsockopt SO_REUSEADDR failed')
		close_socket(server_fd)
		return -1
	}
	if C.setsockopt(server_fd, C.SOL_SOCKET, C.SO_REUSEPORT, &opt, sizeof(opt)) < 0 {
		eprintln(@LOCATION)
		C.perror(c'setsockopt SO_REUSEPORT failed')
		close_socket(server_fd)
		return -1
	}

	addr := if server.family == .ip6 {
		net.new_ip6(u16(server.port), [u8(0), 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]!)
	} else {
		net.new_ip(u16(server.port), [u8(0), 0, 0, 0]!)
	}
	alen := addr.len()
	if C.bind(server_fd, voidptr(&addr), alen) < 0 {
		eprintln(@LOCATION)
		C.perror(c'Bind failed')
		close_socket(server_fd)
		return -1
	}
	if C.listen(server_fd, max_connection_size) < 0 {
		eprintln(@LOCATION)
		C.perror(c'Listen failed')
		close_socket(server_fd)
		return -1
	}
	return server_fd
}

// Function to add a file descriptor to the epoll instance
fn add_fd_to_epoll(epoll_fd int, fd int, events u32) int {
	mut ev := C.epoll_event{
		events: events
	}
	ev.data.fd = fd
	if C.epoll_ctl(epoll_fd, C.EPOLL_CTL_ADD, fd, &ev) == -1 {
		eprintln(@LOCATION)
		C.perror(c'epoll_ctl')
		return -1
	}
	return 0
}

// Function to remove a file descriptor from the epoll instance
fn remove_fd_from_epoll(epoll_fd int, fd int) bool {
	ret := C.epoll_ctl(epoll_fd, C.EPOLL_CTL_DEL, fd, C.NULL)
	if ret == -1 {
		eprintln('ERROR: epoll_ctl(DEL, fd=${fd}) failed with errno=${C.errno}')
		return false
	}
	return true
}

fn handle_accept_loop(epoll_fd int, listen_fd int) {
	for {
		client_fd := C.accept4(listen_fd, C.NULL, C.NULL, C.SOCK_NONBLOCK)
		if client_fd < 0 {
			if C.errno == C.EAGAIN || C.errno == C.EWOULDBLOCK {
				break // No more incoming connections; exit loop.
			}
			eprintln(@LOCATION)
			C.perror(c'Accept failed')
			break
		}
		// Enable TCP_NODELAY for lower latency
		opt := 1
		C.setsockopt(client_fd, C.IPPROTO_TCP, C.TCP_NODELAY, &opt, sizeof(opt))
		// Register client socket with epoll
		if add_fd_to_epoll(epoll_fd, client_fd, u32(C.EPOLLIN | C.EPOLLET)) == -1 {
			close_socket(client_fd)
		}
	}
}

fn handle_client_closure(epoll_fd int, client_fd int) {
	// Never close the listening socket here
	if client_fd == 0 {
		return
	}
	if client_fd <= 0 {
		eprintln('ERROR: Invalid FD=${client_fd} for closure')
		return
	}
	remove_fd_from_epoll(epoll_fd, client_fd)
	close_socket(client_fd)
}

fn process_events(mut server Server, epoll_fd int, listen_fd int) {
	mut events := [max_connection_size]C.epoll_event{}
	mut request_buffer := []u8{len: server.max_request_buffer_size, cap: server.max_request_buffer_size}
	unsafe {
		request_buffer.flags.set(.noslices | .nogrow | .noshrink)
	}
	for {
		num_events := C.epoll_wait(epoll_fd, &events[0], max_connection_size, -1)
		for i := 0; i < num_events; i++ {
			client_fd := unsafe { events[i].data.fd }
			// Accept new connections when the listening socket is readable
			if client_fd == listen_fd {
				handle_accept_loop(epoll_fd, listen_fd)
				continue
			}

			if events[i].events & u32((C.EPOLLHUP | C.EPOLLERR)) != 0 {
				if client_fd == listen_fd {
					eprintln('ERROR: listen fd had HUP/ERR')
					continue
				}
				if client_fd > 0 {
					// Try to send 444 No Response before closing abnormal connection
					C.send(client_fd, status_444_response.data, status_444_response.len,
						C.MSG_NOSIGNAL)
					handle_client_closure(epoll_fd, client_fd)
				} else {
					eprintln('ERROR: Invalid FD from epoll: ${client_fd}')
				}
				continue
			}
			if events[i].events & u32(C.EPOLLIN) != 0 {
				// Read all available data from the socket
				mut total_bytes_read := 0
				mut readed_request_buffer := []u8{cap: server.max_request_buffer_size}

				for {
					bytes_read := C.recv(client_fd, unsafe { &request_buffer[0] }, server.max_request_buffer_size - 1,
						0)
					if bytes_read < 0 {
						if C.errno == C.EAGAIN || C.errno == C.EWOULDBLOCK {
							// No more data available right now
							break
						}
						// Error occurred
						eprintln('ERROR: recv() failed with errno=${C.errno}')
						break
					} else if bytes_read == 0 {
						// Connection closed by client
						break
					}

					// Append the received data to the buffer
					if total_bytes_read + bytes_read > server.max_request_buffer_size {
						// Buffer size exceeded
						break
					}
					unsafe {
						readed_request_buffer.push_many(&request_buffer[0], bytes_read)
					}
					total_bytes_read += bytes_read

					// Check if we've received the complete HTTP request (look for \r\n\r\n)
					if total_bytes_read >= 4 {
						if readed_request_buffer[total_bytes_read - 4] == `\r`
							&& readed_request_buffer[total_bytes_read - 3] == `\n`
							&& readed_request_buffer[total_bytes_read - 2] == `\r`
							&& readed_request_buffer[total_bytes_read - 1] == `\n` {
							break
						}
					}
				}

				if total_bytes_read > 0 {
					// Check if request exceeds buffer size
					if total_bytes_read >= server.max_request_buffer_size - 1 {
						C.send(client_fd, status_413_response.data, status_413_response.len,
							C.MSG_NOSIGNAL)
						handle_client_closure(epoll_fd, client_fd)
						continue
					}
					mut decoded_http_request := decode_http_request(readed_request_buffer) or {
						eprintln('Error decoding request ${err}')
						C.send(client_fd, tiny_bad_request_response.data, tiny_bad_request_response.len,
							C.MSG_NOSIGNAL)
						handle_client_closure(epoll_fd, client_fd)
						continue
					}
					decoded_http_request.client_conn_fd = client_fd
					decoded_http_request.user_data = server.user_data
					response := server.request_handler(decoded_http_request) or {
						eprintln('Error handling request ${err}')
						C.send(client_fd, tiny_bad_request_response.data, tiny_bad_request_response.len,
							C.MSG_NOSIGNAL)
						handle_client_closure(epoll_fd, client_fd)
						continue
					}
					// Send response content (headers/body)
					if response.content.len > 0 {
						mut send_error := false
						mut pos := 0
						for pos < response.content.len {
							sent := C.send(client_fd, unsafe { &response.content[pos] },
								response.content.len - pos, C.MSG_NOSIGNAL)
							if sent <= 0 {
								eprintln('ERROR: send() failed with errno=${C.errno}')
								send_error = true
								break
							}
							pos += sent
						}
						if send_error {
							handle_client_closure(epoll_fd, client_fd)
							continue
						}
					}

					// Send file if present
					if response.file_path != '' {
						fd := C.open(response.file_path.str, C.O_RDONLY)
						if fd == -1 {
							eprintln('ERROR: open file failed')
							handle_client_closure(epoll_fd, client_fd)
							continue
						}
						mut st := C.stat{}
						if C.fstat(fd, &st) != 0 {
							eprintln('ERROR: fstat failed')
							handle_client_closure(epoll_fd, client_fd)
							continue
						}
						mut offset := i64(0)
						mut remaining := i64(st.st_size)
						mut sf_retries := 0
						for remaining > 0 {
							ssize := C.sendfile(client_fd, fd, &offset, usize(remaining))
							if ssize > 0 {
								remaining -= i64(ssize)
								sf_retries = 0
								continue
							}
							errno_val := C.errno
							match errno_val {
								C.EAGAIN, C.EWOULDBLOCK, C.EINTR {
									if sf_retries < 3 {
										sf_retries++
										continue
									}
									eprintln('ERROR: sendfile() transient failure after ${sf_retries} retries (errno=${errno_val})')
								}
								C.EBADF {
									eprintln('ERROR: sendfile() EBADF: input fd or socket not open for required access (errno=${errno_val})')
								}
								C.EFAULT {
									eprintln('ERROR: sendfile() EFAULT: bad address for offset (errno=${errno_val})')
								}
								C.EINVAL {
									eprintln('ERROR: sendfile() EINVAL: invalid descriptor state or non-seekable input (errno=${errno_val})')
								}
								C.EIO {
									eprintln('ERROR: sendfile() EIO: I/O error while reading input file (errno=${errno_val})')
								}
								C.ENOMEM {
									eprintln('ERROR: sendfile() ENOMEM: insufficient kernel memory (errno=${errno_val})')
								}
								C.EOVERFLOW {
									eprintln('ERROR: sendfile() EOVERFLOW: count exceeds file/socket limits (errno=${errno_val})')
								}
								C.ESPIPE {
									eprintln('ERROR: sendfile() ESPIPE: input file not seekable with offset (errno=${errno_val})')
								}
								else {
									eprintln('ERROR: sendfile() failed with errno=${errno_val}')
								}
							}
							handle_client_closure(epoll_fd, client_fd)
							break
						}

						C.close(fd)
					}
					// Leave the connection open; closure is driven by client FIN or errors
				} else if total_bytes_read == 0 {
					// Normal client closure (FIN received)
					handle_client_closure(epoll_fd, client_fd)
				} else if total_bytes_read < 0 && C.errno != C.EAGAIN && C.errno != C.EWOULDBLOCK {
					// Unexpected recv error - send 444 No Response
					C.send(client_fd, status_444_response.data, status_444_response.len,
						C.MSG_NOSIGNAL)
					handle_client_closure(epoll_fd, client_fd)
				}
			}
		}
	}
}

// run starts the server and begins listening for incoming connections.
pub fn (mut server Server) run() ! {
	$if windows {
		eprintln('Windows is not supported yet')
		return
	}
	for i := 0; i < max_thread_pool_size; i++ {
		server.listen_fds[i] = create_server_socket(server)
		if server.listen_fds[i] < 0 {
			return
		}

		server.epoll_fds[i] = C.epoll_create1(0)
		if server.epoll_fds[i] < 0 {
			C.perror(c'epoll_create1 failed')
			close_socket(server.listen_fds[i])
			return
		}

		// Register the listening socket with each worker epoll for distributed accepts (edge-triggered)
		if add_fd_to_epoll(server.epoll_fds[i], server.listen_fds[i], u32(C.EPOLLIN | C.EPOLLET)) == -1 {
			close_socket(server.listen_fds[i])
			close_socket(server.epoll_fds[i])
			return
		}

		server.threads[i] = spawn process_events(mut server, server.epoll_fds[i], server.listen_fds[i])
	}

	println('listening on http://0.0.0.0:${server.port}/')
	// Main thread waits for workers; accepts are handled in worker epoll loops
	for i in 0 .. max_thread_pool_size {
		server.threads[i].wait()
	}
}
